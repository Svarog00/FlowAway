    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   	SavedData   xyhealthcurrentScenemedkitCountquestValues    xSystem.Collections.Generic.List`1[[QuestStages, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   ��?@��?d      ExperementalScene   	      xSystem.Collections.Generic.List`1[[QuestStages, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  QuestStages[]   	                    QuestStages   	   	   	      QuestStages   namestage    	   PowerShield         
   Invisibility            Dash   