    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   	SavedData   xyhealthcurrentScenemedkitCount       �z��� �d      	CityLevel   