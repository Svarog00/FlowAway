    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   	WorldData   xyHealthCurrentSceneMedkitCountQuestValuesItemsAbilityStatuses    wSystem.Collections.Generic.List`1[[QuestStage, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]�System.Collections.Generic.List`1[[System.Boolean, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   ���>r��?d      	CityLevel   	   	   	      wSystem.Collections.Generic.List`1[[QuestStage, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  QuestStage[]   	             ~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  	              �System.Collections.Generic.List`1[[System.Boolean, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  		                    
QuestStage   	
   	   	   	   	          	        
   
QuestStage   	QuestNameStage       Dash      
      SpawnedPlayer      
      MysteriousProblem       
      Invisibility      
      GargoyleFirstMeet    